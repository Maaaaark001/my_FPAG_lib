`define CPOL 0      //clock polarity
`define CPHA 0      //clock phase
`define CLK_FREQ 50_000_000  // input clk frequency
`define SCLK_FREQ  5_000_000  // sclk frequency
`define DATA_WIDTH 8            // a word width
`define CLK_CYCLE 20
